`define INWVAL 24
`define MVAL 5
`define NVAL 4
`define MAXKVAL 6
`define TVPR 0.3
