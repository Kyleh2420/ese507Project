`define OUTWVAL 17
`define DEPTHVAL 48
`define WRENPR 0.01
`define TRPR 0.99
