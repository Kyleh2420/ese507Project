`define INWVAL 24
`define MVAL 5
`define NVAL 4
`define MAXKVAL 2
`define TVPR 0.3
